module adder( a, b, c, q);

input	[3:0]	a,b;
output	[3:0]	q;

assign	q = a + b;

endmodule
